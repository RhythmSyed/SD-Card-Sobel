// $Id: $
// File name:   height_calculator.sv
// Created:     4/14/2018
// Author:      Peiyuan Li
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: calculate the height of the image header
