// $Id: $
// File name:   width_calculator.sv
// Created:     4/14/2018
// Author:      Peiyuan Li
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: calculate the width of the image header.
